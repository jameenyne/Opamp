* spice file for simple amplifier
.include opamp.lib
VDD VDD 0 1.0
VSS VSS 0 -1.0
VS IN 0 0.0
R1 IN NEG 1K
R2 OUT NEG 10K
X1 0 NEG OUT VDD VSS opamp PARAMS: D0=0.034219455569505244 D1=0.04331896697712577 D2=0.04120134893092967 D3=-0.03277415200638261
+    D4=0.015126912454181605 D5=0.016368405175938107 D6=-0.0049206788002917985 D7=-0.023994129007337328 D8=0.003658432372248558
.dc VS -1.0 1.0 0.005
.print dc v(OUT)
.end
